package S_AES_Package;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "S_AES_Seq_Item.svh"
    `include "S_AES_Sequence.svh"
    `include "S_AES_Sequencer.svh"
    `include "S_AES_Driver.svh"
    `include "S_AES_Monitor.svh"
    `include "S_AES_Agent.svh"
    `include "S_AES_Reference_Model.svh"
    `include "S_AES_Scoreboard.svh"
    `include "S_AES_Coverage_Collector.svh"
    `include "S_AES_Env.svh"
    `include "S_AES_Test.sv"

endpackage